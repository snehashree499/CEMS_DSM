** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/Folded Cascode/tb_FolCas_ac.sch
**.subckt tb_FolCas_ac
Vdd v_dd GND 1.8
Vss v_ss GND 0
C1 v_out v_ss 17.98f m=1
Vin v_in v_ss dc 0.8 ac 1
I0 v_dd net1 3u
.save v(v_in)
.save v(v_out)
x1 v_dd net1 v_in v_out v_out v_ss FoldedCascodeOTA
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt

 .lib cornerRES.lib res_typ



.temp 27
.control
option sparse
save all
op
write tb_FolCas_ac.raw
set appendwrite

ac dec 101 1k 1G
write tb_FolCas_ac.raw
plot 20*log10(v_out)

meas ac dcgain MAX vmag(v_out) FROM=10 TO=10k
let f3db = dcgain/sqrt(2)
meas ac fbw WHEN vmag(v_out)=f3db FALL=1
let gainerror=(dcgain-1)/1
print dcgain
print fbw
print gainerror



plot 180/pi*ph(v_out) vs frequency

noise v(v_out) Vin dec 101 1k 100MEG
print onoise_total

.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/Folded Cascode/FoldedCascodeOTA.sym # of pins=6
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/Folded Cascode/FoldedCascodeOTA.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/Folded Cascode/FoldedCascodeOTA.sch
.subckt FoldedCascodeOTA VDD I PLUS MINUS Vout VSS
*.ipin PLUS
*.ipin MINUS
*.opin Vout
*.ipin VDD
*.ipin VSS
*.ipin I
XM1 net2 net4 VDD VDD sg13_lv_pmos w=0.75u l=0.4u ng=1 m=1
XM2 net1 PLUS net2 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM3 net6 MINUS net2 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM14 VSS net9 net6 VSS sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM13 net6 I Vout VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM11 net1 I net7 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM12 VSS net9 net1 VSS sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM9 net8 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM10 net7 net3 net8 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM4 net5 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM5 Vout net3 net5 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM6 net4 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM8 net3 net3 net4 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM7 VSS net9 net3 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM18 net10 I VDD VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM17 VSS net9 net10 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM16 net9 I I VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM15 VSS net9 net9 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
.ends

.GLOBAL GND
.end

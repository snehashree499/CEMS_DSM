** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/IC_Designs_Hrishi/IdealCircuits/IDEAL_DSM_VCCS.sch
**.subckt IDEAL_DSM_VCCS
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75
Vp1 p1 GND dc 0 pulse(0, {vdd}, 5n, 100p, 100p, {per/2-5n}, {per})
Vp2 p2 GND dc {vdd} pulse({vdd}, 0, 0, 100p, 100p, {per/2+5n}, {per})
S1 Vin net1 p1 GND mysw
S2 net4 net2 p2 GND mysw
S3 net1 net3 p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 1p m=1
C1 net4 vo1 6p m=1
S5 vo1 net5 p1 GND mysw
S6 net7 net6 p2 GND mysw
S7 net5 net3 p2 GND mysw
S8 net6 Vcm p1 GND mysw
C2 net5 net6 1p m=1
C3 net7 net8 3p m=1
x2 vcmp Vdd Vss net3 sg13g2_inv_1
Vresb resb GND dc 0 pwl(0, 0, {per/2}, 0, {per/2+100p} {vdd}
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
E1 vo1 GND net4 Vcm -1000
E2 net8 GND net7 Vcm -1000
x3 p1 vcmp net9 GND net8 Comp_Test-3
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.5 per=1u
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 10u 45m uic
plot vcmp vo1
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 vo2 p1 p2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/Comp_Test-3.sym # of pins=5
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/Comp_Test-3.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/Comp_Test-3.sch
.subckt Comp_Test-3 p1 outm outp MINUS PLUS
*.ipin PLUS
*.ipin MINUS
*.ipin p1
*.opin outp
*.opin outm
XMN3 net4 outp outm VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMP5 net4 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP3 outm p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP1 outm outp net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP2 outp outm net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP4 outp p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP6 net3 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XMN4 net3 outm outp VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMN1 net1 PLUS net4 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN2 net1 MINUS net3 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XM7 GND p1 net1 GND sg13_lv_nmos w=4u l=0.18u ng=1 m=1
VDD net2 GND {vdd}
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/IDEAL_DSM/untitled.sch
**.subckt untitled
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75 ac 1
Vp1 p1 GND dc 0 pulse(0, {vdd}, 5n, 100p, 100p, {per/2-5n}, {per})
Vp2 p2 GND dc {vdd} pulse({vdd}, 0, 0, 100p, 100p, {per/2+5n}, {per})
S1 Vin net1 p1 GND mysw
S2 net3 net2 p2 GND mysw
S3 net1 GND p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 410f m=1
C1 net3 vo1 6.49p m=1
Vresb resb GND dc 0 pwl(0, 0, {per/2}, 0, {per/2+100p} {vdd}
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
S5 vo1 net4 p1 GND mysw
S6 net6 net5 p2 GND mysw
S7 net4 GND p2 GND mysw
S8 net5 Vcm p1 GND mysw
C2 net4 net5 54f m=1
C3 net6 vo2 98f m=1
x1 Vcm vo1 net3 STAGE_5tOTA
x2 Vcm vo2 net6 STAGE_5tOTA
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.8 per=1u
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 10n 30u
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 p1 p2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/STAGE_5tOTA.sym # of pins=3
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/STAGE_5tOTA.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/STAGE_5tOTA.sch
.subckt STAGE_5tOTA Plus Vout Minus
*.ipin Minus
*.opin Vout
*.ipin Plus
Vdd v_dd GND 1.8
Vss v_ss GND 0
I0 v_dd net1 3u
x1 v_dd net1 Vout Plus Minus v_ss 5-T_OTA
.ends


* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/5-T_OTA/5-T_OTA.sym # of pins=6
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/5-T_OTA/5-T_OTA.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/5-T_OTA/5-T_OTA.sch
.subckt 5-T_OTA VDD Ibias Vout PLUS MINUS Vss
*.ipin MINUS
*.ipin PLUS
*.ipin VDD
*.ipin Ibias
*.ipin Vss
*.opin Vout
XM10 Vout net1 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM11 net1 net1 VDD VDD sg13_lv_pmos w=0.4u l=0.375u ng=1 m=1
XM12 net2 PLUS net1 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM13 net2 MINUS Vout Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM14 Vss net4 net2 Vss sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM15 net3 VDD VDD Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM16 Vss net4 net3 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM17 net4 VDD Ibias Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM18 Vss net4 net4 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/tb_A_comp.sch
**.subckt tb_A_comp
Vdiff PLUS MINUS {vdiff}
Vmid MINUS GND {vdd/2}
VDD3 p1 GND dc 0 pulse(0, {vdd}, 1n, 50p, 50p, {per/2-1n}, {per})
x1 p1 outm outp MINUS PLUS A_comp-2
**** begin user architecture code


.param temp=27 per=20n vdd=1.5 per=1u vdiff=1m
.option method=gear reltol=1e-5

.control
save all
tran 10p 4n
alterparam vdiff=100m
reset
tran 10p 4n
plot p1 tran1.outm tran1.outp
plot p1 tran2.outm tran2.outp
.endc


 .lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/A_comp-2.sym # of pins=5
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/A_comp-2.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Sneha/A_comp-2.sch
.subckt A_comp-2 p1 outm outp MINUS PLUS
*.opin outp
*.ipin PLUS
*.ipin MINUS
*.ipin p1
*.opin outm
XMN3 net4 outp outm VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMP5 net3 net2 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP1 outm outp net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP2 outp outm net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP6 net1 net2 net2 net2 sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XMN4 net5 outm outp VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMN1 GND net3 net4 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN2 GND net1 net5 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN5 net8 outp outm VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMP7 net8 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP8 outm p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP9 outm outp net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP10 outp outm net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP11 outp p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP12 net7 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XMN6 net7 outm outp VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMN7 net6 PLUS net8 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN8 net6 MINUS net7 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XM7 GND p1 net6 GND sg13_lv_nmos w=4u l=0.18u ng=1 m=1
VDD1 net2 GND {vdd}
.ends

.GLOBAL GND
.end

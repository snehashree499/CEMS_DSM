** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/IC_Designs_Hrishi/RealCircuits/5-T_OTA/tb_5-T_OTA_tran-1.sch
**.subckt tb_5-T_OTA_tran-1
Vdd v_dd GND 1.5
Vss v_ss GND 0
C1 v_out v_ss 0.47p m=1
Vin v_in v_ss dc 0.8 ac 1
I0 v_dd net1 0.8u
.save v(v_in)
.save v(v_out)
x1 v_dd net1 v_out v_in v_out v_ss 5-T_OTA
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt

 .lib cornerRES.lib res_typ



.temp 27
.ic v(v_vout)=0
.control

tran 0.005u 15u uic
plot v_out

let tstart=0
let vout_limit=0.8*0.99
meas tran tcross WHEN v(v_out)=vout_limit

let tsettle=tcross-tstart
print tsettle

.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/5-T_OTA/5-T_OTA.sym # of pins=6
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/5-T_OTA/5-T_OTA.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/5-T_OTA/5-T_OTA.sch
.subckt 5-T_OTA VDD Ibias Vout PLUS MINUS Vss
*.ipin MINUS
*.ipin PLUS
*.ipin VDD
*.ipin Ibias
*.ipin Vss
*.opin Vout
XM10 Vout net1 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM11 net1 net1 VDD VDD sg13_lv_pmos w=0.4u l=0.375u ng=1 m=1
XM12 net2 PLUS net1 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM13 net2 MINUS Vout Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM14 Vss net4 net2 Vss sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM15 net3 VDD VDD Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM16 Vss net4 net3 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM17 net4 VDD Ibias Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM18 Vss net4 net4 Vss sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
.ends

.GLOBAL GND
.end

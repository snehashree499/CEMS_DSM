** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/IC_Designs_Hrishi/RealCircuits/RealSwitchCap_5-T.sch
**.subckt RealSwitchCap_5-T
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75 ac 1
S1 Vin net1 p1 GND mysw
S2 net3 net2 p2 GND mysw
S3 net1 GND p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 0.3p m=1
C1 net3 vo1 2p m=1
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
S5 vo1 net4 p1 GND mysw
S6 net7 net5 p2 GND mysw
S7 net4 GND p2 GND mysw
S8 net5 Vcm p1 GND mysw
C2 net4 net5 0.2p m=1
C3 net7 vo2 0.7p m=1
x1 net3 vo1 Vcm STAGE
x2 net7 vo2 net6 STAGE
Vp1 p1 GND dc 0 pulse(0, {vdd}, 0, 100n, 100n, 2u, 4.5u)
Vp2 p2 GND dc 0 pulse(0, {vdd}, 2.25u, 100n, 100n, 2u, 4.5u)
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.5
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 10n 30u uic
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 p1 p2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/DSM/Designs_Hrishi/STAGE.sym # of pins=3
** sym_path: /foss/designs/DSM/Designs_Hrishi/STAGE.sym
** sch_path: /foss/designs/DSM/Designs_Hrishi/STAGE.sch
.subckt STAGE Plus Vout Minus
*.ipin Minus
*.opin Vout
*.ipin Plus
Vdd v_dd GND 1.8
Vss v_ss GND 0
I0 v_dd net1 3u
*  x1 -  FoldedCascodeOTA  IS MISSING !!!!
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/tb_idsm2.sch
**.subckt tb_idsm2
Vin vin GND dc {vin}
Vssa vssa GND dc 0
Vres res GND dc {vdd} pwl(0, {vdd}, {per/2}, {vdd}, {per/2+25p}, 0)
Vclk clkin GND pulse({vdd}, 0, {per}, 100p, 100p, {0.5*per}, {per})
Vddd VDD GND dc {vdd}
Vssd VSS GND dc 0
Vdda vdda GND dc {vdd}
Vlo vlo GND dc {vlo}
Vhi vhi GND dc {vhi}
C1 dout GND 50f m=1
x1 vhi vlo vdda vssa vin dout res clkin template_idsm2
**** begin user architecture code


.param temp=27 per=20n N=110
.param vlo=0.3 vhi=0.9 vdd=1.2 vin=0.6
.option method=gear reltol=1e-5
.ic v(x1.x3.out1p)=0
.tran 100p {per*N} uic
.meas tran iavg_ana AVG i(Vdda)
.meas tran iavg_dig AVG i(Vddd)

.control
set wr_singlescale
set wr_vecnames
option numdgt = 3
let index = 1
foreach vin_val 0.35 0.4 0.45 0.5 0.55 0.6 0.65 0.7 0.75 0.8 0.85
  alterparam vin = $vin_val
  reset
  run
  set file = {tb_idsm2_}{$&index}{.txt}
  wrdata $file x1.vout1 x1.vout2 dout x1.p1 x1.p2
  destroy $curplot
  let index = index + 1
end
.endc


 .lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.inc /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sym # of pins=8
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sch
.subckt template_idsm2 vhi vlo vdda vssa vin dout res clkin
*.ipin clkin
*.ipin res
*.ipin vin
*.opin dout
*.ipin vssa
*.ipin vdda
*.ipin vlo
*.ipin vhi
*  x4 -  template_clkgen  IS MISSING !!!!
*  x1 -  template_stage  IS MISSING !!!!
*  x2 -  template_stage  IS MISSING !!!!
*  x3 -  template_comp  IS MISSING !!!!
* noconn #net3
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

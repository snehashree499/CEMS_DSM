** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Real_DSM_Design.sch
**.subckt Real_DSM_Design
Vcm Vcm GND dc {vdd/2}
Vin Vin GND SIN(0.7 1.4 80 0 0 0)
S1 Vin net1 p1 GND mysw
S2 net4 net2 p2 GND mysw
S3 net1 net3 p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 0.3p m=1
C1 net4 vo1 2p m=1
S5 vo1 net5 p2 GND mysw
S6 net7 net6 p1 GND mysw
S7 net5 net3 p1 GND mysw
S8 net6 Vcm p2 GND mysw
C2 net5 net6 0.2p m=1
C3 net7 vo2 0.7p m=1
x2 vcmp Vdd Vss net3 sg13g2_inv_1
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
Vp1 p1 GND dc 0 pulse(0, {vdd}, 0, 100n, 100n, 2u, 4.5u)
Vp2 p2 GND dc 0 pulse(0, {vdd}, 2.25u, 100n, 100n, 2u, 4.5u)
x3 Vcm vo1 net4 VCCS_FolCas
x4 Vcm vo2 net7 VCCS_FolCas
x1 p1 GND vcmp GND vo2 A_comp-2
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.5

.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
reset

run
tran 1u 20m

plot vcmp

set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vcmp p1 p2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/VCCS_FolCas.sym # of pins=3
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/VCCS_FolCas.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/VCCS_FolCas.sch
.subckt VCCS_FolCas Plus Vout Minus
*.ipin Minus
*.opin Vout
*.ipin Plus
Vdd v_dd GND 1.5
Vss v_ss GND 0
I0 v_dd net1 0.8u
x1 v_dd net1 Plus Minus Vout v_ss FoldedCascodeOTA
.ends


* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Comparator_design_Sneha/A_comp-2.sym # of pins=5
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Comparator_design_Sneha/A_comp-2.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Comparator_design_Sneha/A_comp-2.sch
.subckt A_comp-2 p1 outm outp MINUS PLUS
*.opin outp
*.ipin PLUS
*.ipin MINUS
*.ipin p1
*.opin outm
XMN3 net4 outp outm VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMP5 net3 net2 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP1 outm outp net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP2 outp outm net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP6 net1 net2 net2 net2 sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XMN4 net5 outm outp VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMN1 GND net3 net4 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN2 GND net1 net5 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN5 net8 outp outm VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMP7 net8 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP8 outm p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP9 outm outp net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP10 outp outm net2 net2 sg13_lv_pmos w=2u l=0.18u ng=1 m=1
XMP11 outp p1 net2 net2 sg13_lv_pmos w=0.5u l=0.18u ng=1 m=1
XMP12 net7 p1 net2 net2 sg13_lv_pmos w=0.5u l=0.15u ng=1 m=1
XMN6 net7 outm outp VSS sg13_lv_nmos w=1u l=0.18u ng=1 m=1
XMN7 net6 PLUS net8 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XMN8 net6 MINUS net7 VSS sg13_lv_nmos w=2u l=0.18u ng=1 m=1
XM7 GND p1 net6 GND sg13_lv_nmos w=4u l=0.18u ng=1 m=1
VDD1 net2 GND {vdd}
.ends


* expanding   symbol:  FoldedCascodeOTA.sym # of pins=6
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sch
.subckt FoldedCascodeOTA VDD I PLUS MINUS Vout VSS
*.ipin PLUS
*.ipin MINUS
*.opin Vout
*.ipin VDD
*.ipin VSS
*.ipin I
XM1 net2 net4 VDD VDD sg13_lv_pmos w=0.272u l=0.5u ng=1 m=1
XM14 VSS net7 net6 VSS sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM13 net6 I Vout VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM11 net1 I net3 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM12 VSS net7 net1 VSS sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM9 net4 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM4 net5 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM6 net4 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM8 net3 net3 net4 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM5 Vout net3 net5 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM10 net3 net3 net4 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM3 net6 MINUS net2 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM2 net1 PLUS net2 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM7 VSS net7 net3 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM18 net8 I VDD VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM17 VSS net7 net8 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM16 net7 I I VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM15 VSS net7 net7 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/IDEAL_DSM/IDEAL_SwitchCap.sch
**.subckt IDEAL_SwitchCap
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75
Vp1 p1 GND dc 0 pulse(0, {vdd}, 5n, 100p, 100p, {per/2-5n}, {per})
Vp2 p2 GND dc {vdd} pulse({vdd}, 0, 0, 100p, 100p, {per/2+5n}, {per})
S1 Vin net1 p1 GND mysw
S2 net4 net2 p2 GND mysw
S3 net1 net3 p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 1p m=1
C1 net4 vo1 6p m=1
S5 vo1 net5 p1 GND mysw
S6 net7 net6 p2 GND mysw
S7 net5 net3 p2 GND mysw
S8 net6 Vcm p1 GND mysw
C2 net5 net6 1p m=1
C3 net7 vo2 3p m=1
E3 vcmp GND TABLE {V(vo2,0)} = (-0.1mV, 0V) (0.1mV, {vdd})
x1 p1 vcmp net8 net9 resb VDD VSS sg13g2_dfrbp_1
x2 vcmp Vdd Vss net3 sg13g2_inv_1
Vresb resb GND dc 0 pwl(0, 0, {per/2}, 0, {per/2+100p} {vdd}
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
E1 vo1 GND net4 Vcm -1000
E2 vo2 GND net7 Vcm -1000
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd=1.2 per=1u
.model mysw SW vt={vdd/2} ron=10k roff=10gig
.option method=gear reltol=1e-4

.control
save all
tran 10n 65u
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata tb_ideal_idsm2.txt vo1 vo2 p1 p2
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/LoopGain.sch
**.subckt LoopGain
C3 vr1 v_ss 0.47p m=1
I3 v_dd Ib 0.8u
Vtest2 vf1 vr1 dc 0 ac 1
C4 net1 v_ss 0.47p m=1
Itest2 v_ss net3 dc 0 ac 1
Vir2 net1 net3 0
.save i(vir2)
Vif2 net3 net2 0
.save i(vif2)
Vdd v_dd GND 1.5
Vss v_ss GND 0
Vin v_in v_ss dc 0.5
x1 v_dd Ib vr1 vf1 v_in v_ss Telescopic
x3 v_dd Ib net1 net2 v_in v_ss Telescopic
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-15
.control
save all

* Operating Point Analysis
op
remzerovec
write tb-loopgain.raw
set appendwrite

* AC Analysis
ac dec 101 1 100G
remzerovec
write tb-loopgain.raw
set appendwrite

* Middlebrook's Method
let tv=-v(vr1)/v(vf1)
let ti=-i(vir1)/i(vif1)
let tmb=(tv*ti - 1)/(tv + ti + 2)

plot db(tmb) ylabel 'Magnitude - Middlebrook'
plot 180/pi*cphase(tmb) ylabel 'Phase - Middlebrook'




*quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sym # of pins=6
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sch
.subckt Telescopic Vdd Ibias1 Vout Vinm Vinp Vss
*.ipin Vinp
*.opin Vout
*.ipin Vinm
*.ipin Vss
*.ipin Vdd
*.ipin Ibias1
XM19 Vss net7 net1 Vss sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM11 net1 Vinp net2 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM14 net1 Vinm net3 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM20 Vout net5 net4 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM25 net9 net5 net10 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM1 Vss net7 net5 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM2 Vss net7 net8 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM3 net8 Ibias1 Vdd Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM4 net3 Ibias1 Vout Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM5 net2 Ibias1 net9 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM6 net4 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM7 net6 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM8 net5 net5 net6 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM9 net10 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM10 Vss net7 net7 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM12 net7 Ibias1 Ibias1 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
.ends

.GLOBAL GND
.end

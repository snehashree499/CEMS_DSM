** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/RealSwitchCap_using_FolCas_OTA.sch
**.subckt RealSwitchCap_using_FolCas_OTA
Vcm Vcm GND dc {vdd/2}
Vin Vin net7 SIN(0 0.7 80 0 0 0)
S1 Vin net1 p1 GND mysw
S2 net3 net2 p2 GND mysw
S3 net1 GND p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 0.3p m=1
C1 net3 vo1 2.06p m=1
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
S5 vo1 net4 p2 GND mysw
S6 net6 net5 p1 GND mysw
S7 net4 GND p1 GND mysw
S8 net5 Vcm p2 GND mysw
C2 net4 net5 0.2p m=1
C3 net6 vo2 0.7p m=1
x1 Vcm vo1 net3 VCCS_FolCas
Vp1 p1 GND dc 0 pulse(0, {vdd}, 0, 100n, 100n, 2u, 4.5u)
Vp2 p2 GND dc 0 pulse(0, {vdd}, 2.25u, 100n, 100n, 2u, 4.5u)
x2 Vcm vo2 net6 VCCS_FolCas
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.5
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 10n 240u
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 vo2 p1 p2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/VCCS_FolCas.sym # of pins=3
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/VCCS_FolCas.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/VCCS_FolCas.sch
.subckt VCCS_FolCas Plus Vout Minus
*.ipin Minus
*.opin Vout
*.ipin Plus
Vdd v_dd GND 1.8
Vss v_ss GND 0
I0 v_dd net1 3u
x1 v_dd net1 Plus Minus Vout v_ss FoldedCascodeOTA
.ends


* expanding   symbol:  /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/Folded
*+ Cascode/FoldedCascodeOTA.sym # of pins=6
** sym_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sym
** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/IC_Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sch
.subckt FoldedCascodeOTA VDD I PLUS MINUS Vout VSS
*.ipin PLUS
*.ipin MINUS
*.opin Vout
*.ipin VDD
*.ipin VSS
*.ipin I
XM1 net2 net4 VDD VDD sg13_lv_pmos w=0.75u l=0.4u ng=1 m=1
XM2 net1 PLUS net2 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM3 net6 MINUS net2 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM14 VSS net9 net6 VSS sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM13 net6 I Vout VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM11 net1 I net7 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM12 VSS net9 net1 VSS sg13_lv_nmos w=0.26u l=0.6u ng=1 m=1
XM9 net8 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM10 net7 net3 net8 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM4 net5 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM5 Vout net3 net5 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM6 net4 net4 VDD VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM8 net3 net3 net4 VDD sg13_lv_pmos w=0.375u l=0.4u ng=1 m=1
XM7 VSS net9 net3 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM18 net10 I VDD VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM17 VSS net9 net10 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM16 net9 I I VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
XM15 VSS net9 net9 VSS sg13_lv_nmos w=0.13u l=0.6u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/tb_Telescopic_ac.sch
**.subckt tb_Telescopic_ac
Vss v_ss GND 0
Vdd v_dd GND 1.5
Vin v_in v_ss dc 0.7 ac 1
.save v(v_in)
I0 v_dd net1 0.8u
C1 v_out v_ss 0.47p m=1
.save v(v_out)
x1 v_dd net1 v_out v_out v_in v_ss Telescopic
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt

 .lib cornerRES.lib res_typ



.temp 27
.control
option sparse
save all
op
write Telescopic_ac.raw
set appendwrite

ac dec 101 1k 0.1G
write Telescopic_ac.raw
plot 20*log10(v_out)

meas ac dcgain MAX vmag(v_out) FROM=10 TO=10k
let f3db = dcgain/sqrt(2)
meas ac fbw WHEN vmag(v_out)=f3db FALL=1
let gainerror=(dcgain-1)/1
print dcgain
print fbw
print gainerror





plot 180/pi*ph(v_out) vs frequency

noise v(v_out) Vin dec 101 1k 100MEG
print onoise_total

.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sym # of pins=6
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Telescopic/Telescopic.sch
.subckt Telescopic Vdd Ibias1 Vout Vinm Vinp Vss
*.ipin Vinp
*.opin Vout
*.ipin Vinm
*.ipin Vss
*.ipin Vdd
*.ipin Ibias1
XM19 Vss net7 net1 Vss sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM11 net1 Vinp net2 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM14 net1 Vinm net3 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM20 Vout net5 net4 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM25 net9 net5 net10 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM1 Vss net7 net5 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM2 Vss net7 net8 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM3 net8 Ibias1 Vdd Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM4 net3 Ibias1 Vout Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM5 net2 Ibias1 net9 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM6 net4 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM7 net6 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM8 net5 net5 net6 Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM9 net10 net6 Vdd Vdd sg13_lv_pmos w=0.16u l=0.5u ng=1 m=1
XM10 Vss net7 net7 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM12 net7 Ibias1 Ibias1 Vss sg13_lv_nmos w=0.15u l=2u ng=1 m=1
.ends

.GLOBAL GND
.end

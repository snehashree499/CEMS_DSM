** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/IC_Designs_Hrishi/IdealCircuits/IdealSwitchCap_VCCS.sch
**.subckt IdealSwitchCap_VCCS
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75 ac 1
S1 Vin net1 p1 GND mysw
S2 net3 net2 p2 GND mysw
S3 net1 GND p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 0.3p m=1
C1 net3 vo1 2.06p m=1
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
S5 vo1 net4 p1 GND mysw
S6 net6 net5 p2 GND mysw
S7 net4 GND p2 GND mysw
S8 net5 Vcm p1 GND mysw
C2 net4 net5 0.2p m=1
C3 net6 vo2 0.7p m=1
G1 GND vo1 Vcm net3 10e-06
G2 GND vo2 Vcm net6 10e-06
Vp1 p1 GND dc 0 pulse(0, {vdd}, 0, 100n, 100n, 2u, 4.5u)
Vp2 p2 GND dc 0 pulse(0, {vdd}, 2.25u, 100n, 100n, 2u, 4.5u)
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.5
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 40u 40u uic
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 p1 p2
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end

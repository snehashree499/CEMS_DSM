** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/tb_FolCas_tran.sch
**.subckt tb_FolCas_tran
Vdd v_dd GND 1.5
Vss v_ss GND 0
C1 v_out v_ss 0.47p m=1
Vin v_in v_ss dc 0.5 ac 1
I0 v_dd net1 0.8u
.save v(v_in)
.save v(v_out)
x1 v_dd net1 v_in v_out v_out v_ss FoldedCascodeOTA
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt

 .lib cornerRES.lib res_typ



.temp 27
.ic v(v_vout)=0
.control

tran 0.005u 15u uic
plot v_out

let tstart=0
let vout_limit = 0.5*0.99
meas tran tcross WHEN v(v_out)=vout_limit

let tsettle=tcross-tstart
print tsettle

.endc


**** end user architecture code
**.ends

* expanding   symbol:  FoldedCascodeOTA.sym # of pins=6
** sym_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sym
** sch_path: /foss/designs/CEMS_DSM/DSM/Schematics/Designs_Hrishi/RealCircuits/Folded Cascode/FoldedCascodeOTA.sch
.subckt FoldedCascodeOTA VDD I PLUS MINUS Vout VSS
*.ipin PLUS
*.ipin MINUS
*.opin Vout
*.ipin VDD
*.ipin VSS
*.ipin I
XM1 net2 net4 VDD VDD sg13_lv_pmos w=0.272u l=0.5u ng=1 m=1
XM14 VSS net7 net6 VSS sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM13 net6 I Vout VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM11 net1 I net3 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM12 VSS net7 net1 VSS sg13_lv_nmos w=0.3u l=2u ng=1 m=1
XM9 net4 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM4 net5 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM6 net4 net4 VDD VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM8 net3 net3 net4 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM5 Vout net3 net5 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM10 net3 net3 net4 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM3 net6 MINUS net2 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM2 net1 PLUS net2 VDD sg13_lv_pmos w=0.136u l=0.5u ng=1 m=1
XM7 VSS net7 net3 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM18 net8 I VDD VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM17 VSS net7 net8 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM16 net7 I I VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
XM15 VSS net7 net7 VSS sg13_lv_nmos w=0.15u l=2u ng=1 m=1
.ends

.GLOBAL GND
.end

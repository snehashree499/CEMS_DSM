** sch_path: /foss/designs/SecondOrder_SingleBit_DSM/DSM/Designs_Hrishi/IDEAL_DSM/IdealSwitchCapacitor.sch
**.subckt IdealSwitchCapacitor
Vcm Vcm GND dc {vdd/2}
Vin Vin GND dc 0.75 ac 1
Vp1 p1 GND dc 0 pulse(0, {vdd}, 5n, 100p, 100p, {per/2-5n}, {per})
Vp2 p2 GND dc {vdd} pulse({vdd}, 0, 0, 100p, 100p, {per/2+5n}, {per})
S1 Vin net1 p1 GND mysw
S2 net3 net2 p2 GND mysw
S3 net1 GND p2 GND mysw
S4 net2 Vcm p1 GND mysw
C7 net1 net2 410f m=1
C1 net3 vo1 6.49p m=1
Vresb resb GND dc 0 pwl(0, 0, {per/2}, 0, {per/2+100p} {vdd}
Vsup VDD GND dc {vdd}
Vss VSS GND dc 0
S5 vo1 net4 p1 GND mysw
S6 net6 net5 p2 GND mysw
S7 net4 GND p2 GND mysw
S8 net5 Vcm p1 GND mysw
C2 net4 net5 54f m=1
C3 net6 vo2 98f m=1
E2 vo1 GND net3 Vcm -1000
E1 vo2 GND net6 Vcm -1000
**** begin user architecture code

.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.inc /foss/pdks/sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27 vdd = 1.8 per=1u
.model mysw SW vt={vdd/2} ron=0.1
.option method=gear reltol=1e-4

.control
save all
run
tran 10n 30u
plot vo1 vo2
set wr_singlescale
set wr_vecnames
wrdata IDEAL_SwitchCap.txt vo1 p1 p2
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end
